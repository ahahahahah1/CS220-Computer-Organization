module and_operator(r0, r1, r2);
input[31:0] r1, r2;
output[31:0] r0;

assign r0 = r1 & r2;

endmodule
`include "./bgt.v"
module bgt_tb();
    reg [31:0] r0, r1, imm, pc;
    wire [31:0] pc_next;

    bgt uut(.r0(r0), .r1(r1), .imm(imm), .pc(pc), .pc_next(pc_next));

    initial begin
        r0 = 32'b0101_0000_0000_0000_0000_0000_0000_0000;
        r1 = 32'b0010_0000_0000_0000_0000_0000_0000_0000;
        imm = 32'b0000_0000_0000_0000_0000_0000_0000_0010;
        pc = 1;
        #10
        r0 = 32'b0000_0010_0000_0000_0000_0000_0000_0000;
        r1 = 32'b0100_0100_0001_0101_0001_0100_0000_0000;
        pc = pc_next;
        #10
        r0 = 32'b0010_0000_0000_0000_0000_0000_0000_0000;
        r1 = 32'b1111_1010_0000_0010_0001_0100_0000_0000;
        pc = pc_next;
        #10
        r0 = 32'b0000_0000_0000_0000_0000_0010_0000_0010;
        r1 = 32'b1111_1111_1111_1111_1111_1111_1111_1111;
        pc = pc_next;
        #10
        r0 = 32'b1110_0000_0110_0101_1001_0000_0100_0000;
        r1 = 32'b1010_0000_0010_0010_0100_0100_0110_0010;
        pc = pc_next;
        #10
        r0 = 32'b1010_1001_0100_0000_0100_0001_0000_0000;
        r1 = 32'b0000_0000_1000_0000_0000_0000_0000_0000;
        pc = pc_next;
    end

    initial begin
        $monitor("r0 = %b\nr1 = %b\npc= %b\npc_next = %b\n", r0, r1, pc, pc_next);
    end
endmodule